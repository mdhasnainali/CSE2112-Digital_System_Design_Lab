module not_gate(in, out); // module_name(inputs, outputs)

// Defining input output and wires
input in;
output out;

// Define circuit functionality
assign out = ~in;
endmodule
